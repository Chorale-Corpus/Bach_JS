BZh91AY&SY�ޝQ �_�Pyg���������`�Ô��������8�]p�B(��D� &�ʛMA��C�� i�T���M4�b1=C ɐ0&F�sL��Lф�hшd�� A��J��C@      sL��Lф�hшd�� @���$%<���S'�z�Q������D�_����̑8I��~���������o�����l���вI섂��}�X�����`�(>��q���ϯ�'�}?G������.���V'��R�X�`,B"p$�� Ҕ��A���X�� �R���č��B,`rJ�� �H���6��X�9�<n�r�\���wP��Oi~���=o�dv��H*�H��1c��-�%�te��b��[x0�az�Tċ��te�����&�T����X$L����H���n�FrHp��\�����±LE	`0��bB7�B�^��5��ک�J�[{l(#K�9�'a�22��fY͙�M��`��j�v,�#��p�
��	�G�Ӥu��n&�p�*:�F�3FŤ��u�f��c�fBk��5��Ji��%���5l5�0�e�:�~�`?��'���`0dx��vB��xf&dx��!=`%�I��N+�4�-3.[s�9	Bm�
�l�Ҧ�mBq�I���ı��#5̓��t�/J���$k�	Wt�X�C����-��k�K�]Jj���e���n5�h��Y�$C�uƢ@���\�γ!�x����;��-@�bc���?�N��N��;{�d ^�<X(! �� _=i�����A�І8�g�ͱcu$�[u�;2A���9�������m"o�[��u�[W���{G'��������0���#[j�?[���ftg�����7�~~�қ6j�X��\D���0h{FRԔ�H������69��º(5� q@m#.��{�S���b���1�������I�Od�0rQ����̍�q��A�ณ�=��&$txb;��q5��d�Ѹ��H��q�|y�¦Jwv��XM)��|����xŸ�}�V�`;�@���ʎޅB�L����K�����B��c�pxr��:Y�^�nf���1Ӝy'ۦP���	48���Lɭ��k�V���9�͚s<�L�Ty���`�|Q�8uVMM;7�����]��G���Cw��O�B1�/���ݩ�<�'a�@�J�M���Y��@US�(�ufo�G�D �AZ�`d��66�P�N���c	:4ٍN�'���y;��V�y"����2l�I���G���xm�]�k���gy��&�w���� �z��L�D2�H*,'O֤]3AM��j���))e��(�(\�\��(Iw,Ir�s2)�!�DQs=�� �G��e)u����9�dVK&�-�MHl�VT��J��卼��o�NF� f�����Z�n�p��(�	�{Trx69�8�c�1ܙ:`�g	�1�U�.0�Q�ٝ�L��Z����5ޑ\�qΰn�08������@�ѱ�w������������9������ĸ�ɔ`�w��;��a&�xs�8ͤ�@P:��������H܁�-�x�܇����.1�gh����:�1`ppET�	���a\Ց!]�FؒE ��Χ��v�)Wa;
z�MH7���9ت/��C�2$t�3��34v�)�$瓒���cr��M6s�·9��>\-����b3�5%4�<5$����G��jŲ[-��)��C�9�n�tX��k�2��Yƣ3����.��I4�8N���cXo;8�<4t4�5��y��Y�89�7���A"��
Pg,��d9�9��H,�cK��C�O9u5�.M��&�\t-M��Z�ˬ`z���Dn�@Dvn{qg>��אv|�;y��f�5:1��q�j�7����5QN`ûdϱ�Lk3T��X�'9<�tx�o)��f��m��'Rpq(�'44f9�.���ܛ�G&�^��,���S��U�o�[m��A�w����������٨H�\���_��}��9�d� �1�2Y$�ȱe���Z�,Y%��RMģ]�ri,���XYWX��

Y"��̃%�ԧ8�
%*MQ�u�b�bN)&%I&���	l�H5�;�3K�VQ�`d����͇U�W�Y�:�����}by_���0$�PKO,��a�Cƙ��/���4�ab�� {0�Jy$�ޏM^�$��sA )���l��#�ȪZ�^3��!m_
핊�*"O1�������4ήs�B�H:�=��?)�����?�}(�jB.!��Xs}�b�.�c�!�Fأ�G��@=w�[���o�pc p�N*#�1�"q��y'8e{��Ʒ|�c�;��R�(%YO��6`x����2#����H�H"*�"� H�Q���@�3B,�����|zX�$;"1b9�Ҙ���%,��%*%�"R�,RIK*,X���De��ks�X��:ƿ���O=O���f� ��ꄂǰȟ�� ��~�W�zA�n&��� �&��A��o�|b���o��ʲ$�c�Em掙~(�[�A��ٷ�9R�E�d����4�Ph�r"x+ݨs����6�;�$�cHH:J�؟��~޽*����<����b� ������P4m}E�l6�Z�9�R${����`|�߄H8���e�3+=�3���g���|MH��#����,c"A�����I�js�,��kR}|�]溽9��8�t�Ǹ�nH�@q�&Iq��x�@[�;KO���<Q�J��\`�ħ]Ԏ>`ѡu7A��f[�	�����,N��0�rnN��}�_�������&�ۀ��� �������=���!���"֚�]DQ~��!)ݪ�L�wWeHw��[��ap�W� qxT��%%,B@bJ<�cϯd��﯅��A�֗�2��_��� �>�|oS�H=��"$45�G�*J=z���p�]£�rE8P��ޝQ